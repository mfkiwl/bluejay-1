        5'h0: rd_data_0 = r_0;
        5'h1: rd_data_0 = r_1;
    