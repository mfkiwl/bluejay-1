module top
(
    input a,
    output logic z,
);
    
always_comb
begin
    case ((a))
    SIZE__WORD:
    begin
        a = b;
    end
    OP__LB:
    begin
        a == c;
        a == c + d;
        y == c + d;
    end
    endcase
end

    hi
    hi
    hi
    hi
    hi

endmodule
